module binding_module();
  
  bind dut_top spi_assertion spi_assertion_bind