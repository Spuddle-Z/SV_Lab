//===================================================================== 
/// Description: 
// the interface of uart
// Designer : wangziyao1@sjtu.edu.cn
// ==================================================================== 

/*
This is only the basic interface, you may change it by your own.
But don't change this signal description.
*/
`timescale 1ns/1ps

interface uart_bus(input logic clk,input logic rst_n);
  // Signal Definition
  // =======================================
  logic tx;
  logic rx;

  // Clocking blocks
  // =======================================
  clocking slv_cb @(posedge clk);
    default input #0.25 output #0.25;
    input tx;
    output rx;
  endclocking

  clocking mnt_cb @(posedge clk);
    default input #0.25 output #0.25;
    input tx, rx;
  endclocking

  // Mod ports
  // =======================================
  modport master(
    output tx,
    input rx, clk, rst_n
  );
  modport slave(
    input clk, rst_n,
    clocking slv_cb
  );
  modport monitor(
    input clk, rst_n,
    clocking mnt_cb
  );
endinterface:uart_bus //uart  