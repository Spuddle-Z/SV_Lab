`define SVA