`timescale 1ns/1ps

module spi_slave (
    // --- SPI 引脚（模式 0，低位先行）
    input  logic        sck,     // SPI 时钟
    input  logic        cs_n,    // SPI 片选
    input  logic        mosi,    // 主设备输出，从设备输入
    output logic        miso,    // 主设备输入，从设备输出

    // --- 系统时钟与复位
    input  logic        clk,     // 系统时钟
    input  logic        rst_n,   // 低有效复位

    // --- 数据与控制接口
    input  logic [31:0] tx_data,
    input  logic        tx_valid,
    output logic        tx_done,

    output logic [31:0] rx_data,
    output logic        rx_done
  );

  // ============================================================================
  // 直接使用SPI引脚信号
  // ============================================================================
  logic sck_synced, cs_n_synced, mosi_synced;
  assign sck_synced  = sck;
  assign cs_n_synced = cs_n;
  assign mosi_synced = mosi;

  // ============================================================================
  // 边沿检测
  // ============================================================================
  logic sck_prev, sample_edge, shift_edge;
  logic cs_n_prev, start_edge, stop_edge;

  always_ff @(posedge clk or negedge rst_n) begin
    if (!rst_n) begin
      sck_prev <= 1'b0;
      cs_n_prev <= 1'b1;
    end else begin
      sck_prev <= sck_synced;
      cs_n_prev <= cs_n_synced;
    end
  end

  assign sample_edge = sck_synced && !sck_prev;
  assign shift_edge = !sck_synced && sck_prev;
  assign start_edge = !cs_n_synced && cs_n_prev;
  assign stop_edge = cs_n_synced && !cs_n_prev;

  // ============================================================================
  // 移位寄存器
  // ============================================================================
  logic [31:0] tx_shift_reg;
  logic tx_en;
  logic [5:0] bit_cnt;

  always_ff @(posedge clk or negedge rst_n) begin
    if (!rst_n) begin
      tx_shift_reg <= 32'b0;
      tx_en <= 1'b0;
      bit_cnt <= 6'd0;
    end else begin
      if (start_edge && tx_valid) begin
        tx_shift_reg <= tx_data;
        tx_en <= 1'b1;
        bit_cnt <= 6'd0;
      end else if (!cs_n_synced && sample_edge) begin
        rx_data <= {mosi_synced, rx_data[31:1]};
      end else if (!cs_n_synced && shift_edge && tx_en) begin
        tx_shift_reg <= {1'b0, tx_shift_reg[31:1]};
        if (bit_cnt == 6'd31) begin
          tx_en <= 1'b0;
        end else begin
          bit_cnt <= bit_cnt + 1'b1;
        end
      end else if (stop_edge) begin
        tx_en <= 1'b0;
        bit_cnt <= 6'd0;
      end
    end
  end

  assign rx_done = stop_edge;
  assign tx_done = stop_edge;
  assign miso = tx_en ? tx_shift_reg[0] : 1'b0;

endmodule

module ctrl_reg (
  // 时钟和复位
  input  logic    clk,
  input  logic    rst_n,
  
  // 总线接口
  input  logic [31:0] spi_rx_data,
  input  logic        spi_rx_done,
  output logic [31:0] spi_tx_data,
  output logic        rx_reg_valid,
  input  logic        spi_tx_done,

  // FIFO接口
  output logic [15:0] tx_fifo_data,
  input  logic        tx_fifo_full,
  output logic        tx_fifo_en,
  input  logic [31:0] rx_fifo_data,
  input  logic        rx_fifo_empty,
  output logic        rx_fifo_en,

  // UART控制信号
  input  logic [3:0]  state,
  output logic [15:0] baud,
  output logic [1:0] control
);
  // ============================================================================
  // 寄存器定义
  // ============================================================================
  logic [1:0] control_reg;
  logic [3:0] state_reg;
  logic [15:0] baud_reg;
  logic [31:0] rx_data_reg;

  // ============================================================================
  // 解析命令
  // ============================================================================
  logic [7:0] command, addr;
  logic [15:0] data;

  assign command = spi_rx_data[31:24];
  assign addr    = spi_rx_data[23:16];
  assign data    = spi_rx_data[15:0];

  typedef enum logic [7:0] {
    CONTROL = 8'h00,
    STATE = 8'h08,
    TX_DATA = 8'h10,
    RX_DATA = 8'h18,
    BAUD = 8'h20
  } addr_t;

  // ============================================================================
  // 控制寄存器写逻辑
  // ============================================================================
  always_ff @(posedge clk or negedge rst_n) begin
    if (!rst_n) begin
      control_reg <= 2'b0;
      state_reg <= 4'b0;
      baud_reg <= 16'b0;
      rx_data_reg <= 32'b0;
      spi_tx_data <= 32'b0;
      rx_reg_valid <= 1'b0;
      tx_fifo_en <= 1'b0;
      rx_fifo_en <= 1'b0;
    end else begin // 处理接收到的数据
      tx_fifo_en <= 1'b0;
      rx_fifo_en <= 1'b0;
      if (spi_tx_done)
        rx_reg_valid <= 1'b0;
      if (spi_rx_done) begin
        case (command)
          8'h00: begin
            case (addr)
              CONTROL: control_reg <= data[1:0];
              TX_DATA: begin
                tx_fifo_data <= data;
                tx_fifo_en <= 1'b1;
              end
              BAUD: baud_reg <= data;
            endcase
          end
          8'h01: begin
            rx_reg_valid <= 1'b1;
            case (addr)
              CONTROL: spi_tx_data <= {30'b0, control_reg};
              STATE: spi_tx_data <= {28'b0, state_reg};
              RX_DATA: begin
                spi_tx_data <= rx_data_reg;
                rx_fifo_en <= 1'b1;
              end
              BAUD: spi_tx_data <= {16'b0, baud_reg};
            endcase
          end
        endcase
      end
    end
  end

  // ============================================================================
  // RX_FIFO接收
  // ============================================================================
  always_ff @(posedge clk or negedge rst_n) begin
    if (!rst_n) begin
      rx_data_reg <= 32'b0;
    end else if (rx_fifo_en) begin
      rx_data_reg <= rx_fifo_empty ? 32'h0 : rx_fifo_data;
    end
  end

  // ============================================================================
  // 输出信号赋值
  // ============================================================================
  assign control = control_reg;
  assign baud = baud_reg;

endmodule

module spi_ctl (
  input  logic        clk,
  input  logic        rst_n,

  // SPI引脚
  input  logic        sck,      // SPI时钟
  input  logic        cs_n,     // SPI片选
  input  logic        mosi,     // 主设备输出，从设备输入
  output logic        miso,     // 主设备输入，从设备输出

  // TX FIFO接口
  output logic [15:0] tx_fifo_data,
  input  logic        tx_fifo_full,
  output logic        tx_fifo_en,

  // RX FIFO接口
  input  logic [31:0] rx_fifo_data,
  input  logic        rx_fifo_empty,
  output logic        rx_fifo_en,
  
  // UART控制信号
  input  logic [3:0]  state,
  output logic [1:0]  control,
  output logic [15:0] baud
);

  // ============================================================================
  // 信号定义
  // ============================================================================
  // SPI与控制寄存器接口
  logic [31:0] spi_rx_data;
  logic        spi_rx_done;
  logic [31:0] spi_tx_data;
  logic        rx_reg_valid;
  logic        spi_tx_done;

  // ============================================================================
  // DUT实例化
  // ============================================================================
  spi_slave spi_slave_inst (
    .sck(sck),
    .cs_n(cs_n),
    .mosi(mosi),
    .miso(miso),

    .clk(clk),
    .rst_n(rst_n),

    .rx_data(spi_rx_data),
    .rx_done(spi_rx_done),
    .tx_data(spi_tx_data),
    .tx_valid(rx_reg_valid),
    .tx_done(spi_tx_done)
  );

  ctrl_reg dut (
    .clk(clk),
    .rst_n(rst_n),

    .spi_rx_data(spi_rx_data),
    .spi_rx_done(spi_rx_done),
    .spi_tx_data(spi_tx_data),
    .rx_reg_valid(rx_reg_valid),
    .spi_tx_done(spi_tx_done),

    .tx_fifo_data(tx_fifo_data),
    .tx_fifo_full(tx_fifo_full),
    .tx_fifo_en(tx_fifo_en),
    .rx_fifo_data(rx_fifo_data),
    .rx_fifo_empty(rx_fifo_empty),
    .rx_fifo_en(rx_fifo_en),

    .state(state),
    .control(control),
    .baud(baud)
  );

endmodule